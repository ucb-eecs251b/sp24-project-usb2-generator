* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDM-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
M0 VGND A Y VNB nfet_01v8 w=0.65u l=0.15u
M1 VPWR A Y VPB pfet_01v8_hvt w=1u l=0.15u
M2 Y A VGND VNB nfet_01v8 w=0.65u l=0.15u
M3 Y A VGND VNB nfet_01v8 w=0.65u l=0.15u
M4 VPWR A Y VPB pfet_01v8_hvt w=1u l=0.15u
M5 Y A VPWR VPB pfet_01v8_hvt w=1u l=0.15u
M6 Y A VPWR VPB pfet_01v8_hvt w=1u l=0.15u
M7 Y A VPWR VPB pfet_01v8_hvt w=1u l=0.15u
M8 Y A VPWR VPB pfet_01v8_hvt w=1u l=0.15u
M9 VPWR A Y VPB pfet_01v8_hvt w=1u l=0.15u
M10 VGND A Y VNB nfet_01v8 w=0.65u l=0.15u
M11 Y A VGND VNB nfet_01v8 w=0.65u l=0.15u
M12 Y A VGND VNB nfet_01v8 w=0.65u l=0.15u
M13 VGND A Y VNB nfet_01v8 w=0.65u l=0.15u
M14 VGND A Y VNB nfet_01v8 w=0.65u l=0.15u
M15 VPWR A Y VPB pfet_01v8_hvt w=1u l=0.15u
.ends