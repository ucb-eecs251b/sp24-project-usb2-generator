/scratch/eecs251b-aaz/sp24-project-usb2-generator/build copy/tech-sky130-cache/sky130_ef_io.lef