===================
Spice In Log File
===================
Parameter file: /tmp/spiceInPw63957
Import Parameters:
	Netlist file name: /home/ff/eecs251b/sky130/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
	Output library name: test
	Output View Type: schematic
	Schematic view name: schematic
	Netlist view name: netlist_tmp
	Reference Library List: sky130_fd_pr_main test 
	Top cell: top
	Device-mapping not enabled.
	Master Cell for Ground: gnd
	Schematic Generation parameter file: /tmp/schOpts_spiceInPw63957
	Simulator: spectre
	Output Simulator: spectre
	paramCaseValue: default
	Language: SPICE
Total number of files: 1.

Netlist File: /home/ff/eecs251b/sky130/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice.
Total number of Subckts: 437.

********
Created test.sky130_fd_sc_hd__a2bb2o_1:netlist_tmp
	Created net A1_N.
	Created term A1_N.
	Created net A2_N.
	Created term A2_N.
	Created net B1.
	Created term B1.
	Created net B2.
	Created term B2.
	Created net VGND.
	Created term VGND.
	Created net VNB.
	Created term VNB.
	Created net VPB.
	Created term VPB.
	Created net VPWR.
	Created term VPWR.
	Created net X.
	Created term X.

	Total number of Insts: 12.

	Inst: X0
		Created net 'a_489_413#'.
		Found net 'B2'.
		Found net 'VPWR'.
		Found net 'VPB'.

		Master Cell: 'sky130_fd_pr__pfet_01v8_hvt'.
		Did not find 'sky130_fd_pr_main.sky130_fd_pr__pfet_01v8_hvt:symbol'.
		Did not find test.sky130_fd_pr__pfet_01v8_hvt:schematic.
ERROR (SPICEIN-24): Spice In did not find the symbol view of the master cell 'sky130_fd_pr__pfet_01v8_hvt' of the instance
'X0' in the subcircuit 'sky130_fd_sc_hd__a2bb2o_1'. Specify the reference library that has the symbol
view of the master cell, or use device-mapping to map 'sky130_fd_pr__pfet_01v8_hvt' to a different cell.
Some device mapping file examples for commonly used components while importing
a spice netlist include: 
devselect := resistor res
devselect := capacitor cap
devselect := inductor ind
devselect := mutual_inductor mind
Search 'SPICEIN-24' in Cadence Help for more information.
INFO (SPICEIN-56): Spice In failed to import the netlist file '/home/ff/eecs251b/sky130/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice'. You may like to read the log
file '/scratch/eecs251b-aaz/sp24-project-usb2-generator/cadence/sky130_fd_sc_hd__lpflow_inputisolatch_1.spice' for details.
